module traffic_light_tb;

reg clk;
reg reset;
wire red;
wire yellow;
wire green;

traffic_light UUT (
    .clk(clk),
    .reset(reset),
    .red(red),
    .yellow(yellow),
    .green(green)
);

always #5 clk = ~clk;

initial
begin
    clk = 0;
    reset = 1;

    #10 reset = 0;

    #100 $stop;
end

endmodule

